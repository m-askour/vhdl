library library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nom is 
    port (signaux);
end  nom;

architecture STRUCTURE_DE_BASE of nom is

end STRUCTURE_DE_BASE;